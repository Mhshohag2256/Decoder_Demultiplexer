library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Shohag_3to8Decoder_test is
Port ( 	Shohag_IN : in STD_LOGIC_VECTOR (2 downto 0);
			Shohag_OUT : out STD_LOGIC_VECTOR (7 downto 0));
end Shohag_3to8Decoder_test;

architecture arch of Shohag_3to8Decoder_test is
	begin
	
			with Shohag_IN select
			Shohag_OUT<="00000001" when "000",
				"00000010" when "001",
				"00000100" when "010",
				"00001000" when "011",
				"00010000" when "100",
				"00100000" when "101",
				"01000000" when "110",
				"10000000" when "111",
				"00000000" when others;
end arch;
